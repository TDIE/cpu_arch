//This package contains everything to run the UVM base test for the cpu
//Author: Tom Diederen
//December 2023
//Part of Rudimentary Processor Design Project: https://github.com/TDIE/cpu_arch

package base_test_pkg;
    import uvm_pkg::*;
    import cpu_agent_pkg::*;
    import cpu_env_pkg::*;
    `include "base_test.svh"
    //`include "cpu_bus_seq.svh"
endpackage: base_test_pkg
