//This package contains everything related to the cpu_agent
//Author: Tom Diederen
//December 2023
//Part of Rudimentary Processor Design Project: https://github.com/TDIE/cpu_arch

package cpu_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "cpu_agent.svh"
    // `include "cpu_monitor.svh"
    // `include "cpu_driver.svh"
    // `include "cpu_mon_bus_seq_item.svh"
    // `include "cpu_drv_bus_seq_item.svh"
    // `incluce "cpu_agent_config"
endpackage: cpu_agent_pkg