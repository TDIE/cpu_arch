//This package contains everything related to the cpu_env
//Author: Tom Diederen
//December 2023
//Part of Rudimentary Processor Design Project: https://github.com/TDIE/cpu_arch

package cpu_env_pkg;
    import uvm_pkg::*;
    import cpu_agent_pkg::*;
    `include "uvm_macros.svh"
    `include "cpu_env.svh"
    //`include "scoreboard.svh"
    //`include "coverage_collector.svh"
    //`include "cpu_env_config.svh"
endpackage: cpu_env_pkg